library verilog;
use verilog.vl_types.all;
entity OR16bit_tb is
end OR16bit_tb;
