library verilog;
use verilog.vl_types.all;
entity Testbench is
    generic(
        N               : integer := 16
    );
end Testbench;
