library verilog;
use verilog.vl_types.all;
entity carry_look_ahead_16bit_tb is
end carry_look_ahead_16bit_tb;
