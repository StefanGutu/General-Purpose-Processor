library verilog;
use verilog.vl_types.all;
entity CMP16bit_tb is
end CMP16bit_tb;
