library verilog;
use verilog.vl_types.all;
entity RSR16bit_tb is
end RSR16bit_tb;
