library verilog;
use verilog.vl_types.all;
entity tb_division is
    generic(
        WIDTH           : integer := 16
    );
end tb_division;
