library verilog;
use verilog.vl_types.all;
entity RSL16bit_tb is
end RSL16bit_tb;
