library verilog;
use verilog.vl_types.all;
entity NOT16bit_tb is
end NOT16bit_tb;
