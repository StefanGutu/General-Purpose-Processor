library verilog;
use verilog.vl_types.all;
entity LSL16bit_tb is
end LSL16bit_tb;
