library verilog;
use verilog.vl_types.all;
entity XOR16bit_tb is
end XOR16bit_tb;
