library verilog;
use verilog.vl_types.all;
entity TST16bit_tb is
end TST16bit_tb;
