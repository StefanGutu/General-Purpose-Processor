library verilog;
use verilog.vl_types.all;
entity AND16bit_tb is
end AND16bit_tb;
