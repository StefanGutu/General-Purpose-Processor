library verilog;
use verilog.vl_types.all;
entity DEC16bit_tb is
end DEC16bit_tb;
