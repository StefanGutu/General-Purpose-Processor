library verilog;
use verilog.vl_types.all;
entity MOV16bit_tb is
end MOV16bit_tb;
