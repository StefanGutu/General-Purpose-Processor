library verilog;
use verilog.vl_types.all;
entity tb_FSM16bit is
end tb_FSM16bit;
