library verilog;
use verilog.vl_types.all;
entity INC16bit_tb is
end INC16bit_tb;
