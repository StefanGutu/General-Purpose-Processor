library verilog;
use verilog.vl_types.all;
entity LSR16bit_tb is
end LSR16bit_tb;
