library verilog;
use verilog.vl_types.all;
entity MOD16bit_tb is
end MOD16bit_tb;
