library verilog;
use verilog.vl_types.all;
entity FullSubtractor16bit_tb is
end FullSubtractor16bit_tb;
